<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Associação de Natação de Coimbra" version="11.77730">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Coimbra" name="V Open de Natação Adaptada da Associação de Natação de Coimbra" course="LCM" deadline="2023-11-21" number="1" organizer="ANC" organizer.url="https://www.ancoimbra.pt" reservecount="2" startmethod="1" timing="AUTOMATIC" type="POR.NA" nation="POR" maxentriesathlete="4">
      <AGEDATE value="2023-12-02" type="POR" />
      <POOL name="Centro Olimpico de Piscinas de Coimbra" lanemax="9" />
      <FACILITY city="Coimbra" name="Centro Olimpico de Piscinas de Coimbra" nation="POR" street="Praça Herois do Ultramar - COP" zip="3030-327" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <CONTACT email="geral@ancoimbra.pt" name="Paula Toscano" phone="239855000/917420979" street="Praça Herois do Ultramar - COP" zip="3030-327" />
      <SESSIONS>
        <SESSION date="2023-12-02" daytime="09:30" name="1ª Jornada - 1ª Sessão" number="1" warmupfrom="08:00" warmupuntil="09:15" maxentriesathlete="2">
          <EVENTS>
            <EVENT eventid="1077" daytime="09:30" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15090" agemax="-1" agemin="10" name="Classe S6-S14-Absolutos" handicap="6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="15091" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18090" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="15117" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="15093" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="15094" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="15095" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="15096" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="15097" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="15098" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="15099" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="15100" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="15101" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="15102" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="15103" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="15104" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="15105" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="15106" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="15107" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="15108" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="15109" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="15110" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="15111" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="15112" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="15113" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18091" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18092" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="15118" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="15092" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="15114" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="15115" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="15305" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="15116" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="15119" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1085" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18093" agemax="-1" agemin="10" name="Classe S6-S14-Absolutos" handicap="6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="18094" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18095" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18096" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="18097" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="18098" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="18099" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="18100" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="18101" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="18102" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="18103" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="18104" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="18105" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="18106" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="18107" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="18108" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="18109" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="18110" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="18111" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="18112" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="18113" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="18114" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18115" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18116" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18117" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18118" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18119" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18120" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18121" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18122" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18123" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18124" agemax="-1" agemin="-1" name="Classe S110" />
                <AGEGROUP agegroupid="18125" agemax="-1" agemin="-1" name="Classe S113" />
                <AGEGROUP agegroupid="18126" agemax="-1" agemin="-1" name="Classe S114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1122" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23250" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="23251" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="23252" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="23253" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="23254" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="23255" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="23256" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="23257" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="23258" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="23259" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="23260" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="23261" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="23262" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="23263" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="23264" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="23265" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="23266" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="23267" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="23268" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="23269" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="23270" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="23271" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="23272" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="23273" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="23274" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="23275" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="23276" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="23277" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="23278" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="23279" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="23280" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="23281" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="23282" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="23283" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="23284" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="23285" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="23286" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="23287" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="23288" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="23289" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="23290" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="23291" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="23292" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="23293" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1128" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23294" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="23295" agemax="-1" agemin="8" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="23296" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="23297" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="23298" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="23299" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="23300" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="23301" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="23302" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="23303" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="23304" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="23305" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="23306" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="23307" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="23308" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="23309" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="23310" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="23311" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="23312" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="23313" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="23314" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="23315" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="23316" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="23317" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="23318" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="23319" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="23320" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="23321" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="23322" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="23323" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="23324" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="23325" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="23326" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="23327" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="23328" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="23329" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="23330" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="23331" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="23332" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="23333" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="23334" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="23335" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="23336" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="23337" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1110" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18196" agemax="-1" agemin="10" name="Classe SB4-SB14-Absolutos" handicap="4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="18197" agemax="-1" agemin="10" name="Classe SB15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18198" agemax="-1" agemin="-1" name="Classe SB16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18199" agemax="-1" agemin="-1" name="Classe SB17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="18200" agemax="-1" agemin="10" name="Classe SB21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="18201" agemax="16" agemin="10" name="Classe SB4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="18202" agemax="-1" agemin="17" name="Classe SB4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="18203" agemax="16" agemin="10" name="Classe SB5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="18204" agemax="-1" agemin="17" name="Classe SB5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="18205" agemax="16" agemin="10" name="Classe SB6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="18206" agemax="-1" agemin="17" name="Classe SB6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="18207" agemax="16" agemin="10" name="Classe SB7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="18208" agemax="-1" agemin="17" name="Classe SB7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="18209" agemax="16" agemin="10" name="Classe SB8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="18210" agemax="-1" agemin="17" name="Classe SB8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="18211" agemax="16" agemin="9" name="Classe SB9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="18212" agemax="-1" agemin="17" name="Classe SB9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="18213" agemax="16" agemin="10" name="Classe SB10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="18214" agemax="-1" agemin="17" name="Classe SB10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="18215" agemax="16" agemin="10" name="Classe SB11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="18216" agemax="-1" agemin="17" name="Classe SB11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="18217" agemax="16" agemin="10" name="Classe SB12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="18218" agemax="-1" agemin="17" name="Classe SB12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="18219" agemax="16" agemin="10" name="Classe SB13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="18220" agemax="-1" agemin="17" name="Classe SB13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="18221" agemax="16" agemin="10" name="Classe SB14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18222" agemax="-1" agemin="17" name="Classe SB14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18223" agemax="16" agemin="10" name="Classe SB15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18224" agemax="-1" agemin="17" name="Classe SB15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18225" agemax="16" agemin="10" name="Classe SB16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18226" agemax="-1" agemin="17" name="Classe SB16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18227" agemax="16" agemin="10" name="Classe SB17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18228" agemax="-1" agemin="17" name="Classe SB17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18229" agemax="16" agemin="10" name="Classe SB21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18230" agemax="-1" agemin="17" name="Classe SB21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18231" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="18232" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="18233" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1118" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15179" agemax="-1" agemin="10" name="Classe SB4-SB14-Absolutos" handicap="4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="15180" agemax="-1" agemin="10" name="Classe SB15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18193" agemax="-1" agemin="-1" name="Classe SB16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="15181" agemax="-1" agemin="-1" name="Classe SB17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="15182" agemax="-1" agemin="10" name="Classe SB21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="15183" agemax="16" agemin="10" name="Classe SB4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="15184" agemax="-1" agemin="17" name="Classe SB4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="15185" agemax="16" agemin="10" name="Classe SB5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="15186" agemax="-1" agemin="17" name="Classe SB5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="15187" agemax="16" agemin="10" name="Classe SB6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="15188" agemax="-1" agemin="17" name="Classe SB6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="15189" agemax="16" agemin="10" name="Classe SB7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="15190" agemax="-1" agemin="17" name="Classe SB7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="15191" agemax="16" agemin="10" name="Classe SB8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="15192" agemax="-1" agemin="17" name="Classe SB8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="15193" agemax="16" agemin="9" name="Classe SB9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="15194" agemax="-1" agemin="17" name="Classe SB9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="15195" agemax="16" agemin="10" name="Classe SB10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="15196" agemax="-1" agemin="17" name="Classe SB10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="15197" agemax="16" agemin="10" name="Classe SB11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="15198" agemax="-1" agemin="17" name="Classe SB11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="15199" agemax="16" agemin="10" name="Classe SB12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="15200" agemax="-1" agemin="17" name="Classe SB12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="15201" agemax="16" agemin="10" name="Classe SB13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="15202" agemax="-1" agemin="17" name="Classe SB13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="15203" agemax="16" agemin="10" name="Classe SB14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="15204" agemax="-1" agemin="17" name="Classe SB14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="15205" agemax="16" agemin="10" name="Classe SB15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="15206" agemax="-1" agemin="17" name="Classe SB15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="15207" agemax="16" agemin="10" name="Classe SB16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="15208" agemax="-1" agemin="17" name="Classe SB16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18194" agemax="16" agemin="10" name="Classe SB17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18195" agemax="-1" agemin="17" name="Classe SB17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="15209" agemax="16" agemin="10" name="Classe SB21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="15210" agemax="-1" agemin="17" name="Classe SB21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="15211" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="15212" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="15213" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5931" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18326" agemax="-1" agemin="10" name="Classe S14-Absoluto" handicap="14" />
                <AGEGROUP agegroupid="18327" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absoluto" handicap="15" />
                <AGEGROUP agegroupid="20947" agemax="-1" agemin="10" name="Classe S17-Absoluto" handicap="17" />
                <AGEGROUP agegroupid="18329" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absoluto" handicap="21" />
                <AGEGROUP agegroupid="18330" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18331" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18332" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18333" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18334" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18335" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18336" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18337" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18328" agemax="-1" agemin="10" name="Classe S9-Absoluto" handicap="9" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5916" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18323" agemax="-1" agemin="10" name="Classe S14-Absoluto" handicap="14" />
                <AGEGROUP agegroupid="7728" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absoluto" handicap="15" />
                <AGEGROUP agegroupid="7725" agemax="-1" agemin="10" name="Classe S17-Absoluto" handicap="17" />
                <AGEGROUP agegroupid="7731" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absoluto" handicap="21" />
                <AGEGROUP agegroupid="7726" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="7727" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18324" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18325" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="7729" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="7730" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="7732" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="7733" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="20946" agemax="-1" agemin="10" name="Classe S8" handicap="8" />
                <AGEGROUP agegroupid="20914" agemax="-1" agemin="10" name="Classe S113" handicap="113" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1209" gender="F" number="9" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18409" agemax="-1" agemin="10" name="Classe S8-S14-Absolutos" handicap="8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="18410" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18411" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18412" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="18413" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="18414" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="18415" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="18416" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="18417" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="18418" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="18419" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="18420" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="18421" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="18422" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="18423" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="18424" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="18425" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="18426" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18427" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18428" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18429" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18430" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18431" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18432" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18433" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18434" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18435" agemax="-1" agemin="17" name="Classe S21 (SDown)-Senior" handicap="21" />
                <AGEGROUP agegroupid="18436" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="18437" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="18438" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1201" gender="M" number="10" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7821" agemax="-1" agemin="10" name="Classe S8-S14-Absolutos" handicap="8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="7832" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="15224" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18406" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="7831" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="7825" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="1204" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="7826" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="1205" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="7827" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="1972" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="7828" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="1973" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="7829" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="3971" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="7830" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="1206" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="7822" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="1207" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="7823" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="6013" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="15225" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="6258" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18407" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18408" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="7824" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="1974" agemax="-1" agemin="17" name="Classe S21 (SDown)-Senior" handicap="21" />
                <AGEGROUP agegroupid="3257" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="6259" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="15223" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5946" gender="F" number="11" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18234" agemax="-1" agemin="10" name="Classe S14-Absoluto" handicap="14" />
                <AGEGROUP agegroupid="7674" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absoluto" handicap="15" />
                <AGEGROUP agegroupid="7671" agemax="-1" agemin="10" name="Classe S17-Absoluto" handicap="17" />
                <AGEGROUP agegroupid="7677" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absoluto" handicap="21" />
                <AGEGROUP agegroupid="7672" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="7673" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18235" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18236" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="7675" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="7676" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="7678" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="7679" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="15253" agemax="-1" agemin="17" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5957" gender="M" number="12" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18237" agemax="-1" agemin="10" name="Classe S14-Absoluto" handicap="14" />
                <AGEGROUP agegroupid="18238" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absoluto" handicap="15" />
                <AGEGROUP agegroupid="18239" agemax="-1" agemin="10" name="Classe S17-Absoluto" handicap="17" />
                <AGEGROUP agegroupid="18240" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absoluto" handicap="21" />
                <AGEGROUP agegroupid="18241" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18242" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18243" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18244" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18245" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18246" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18247" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18248" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18249" agemax="-1" agemin="17" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7320" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18442" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="18443" agemax="-1" agemin="8" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18444" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18445" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="18446" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="18447" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="18448" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="18449" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="18450" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="18451" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="18452" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="18453" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="18454" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="18455" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="18456" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="18457" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="18458" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="18459" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="18460" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="18461" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="18462" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="18463" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="18464" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="18465" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="18466" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="18467" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="18468" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="18469" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="18470" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="18471" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="18472" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="18473" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18474" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18475" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18476" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18477" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18478" agemax="-1" agemin="17" name="Classe S16-Senior" handicap="16" />
                <AGEGROUP agegroupid="18479" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18480" agemax="-1" agemin="17" name="Classe S17-Senior" handicap="17" />
                <AGEGROUP agegroupid="18481" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18482" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18483" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="18484" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="18485" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="7322" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="11112" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="7977" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18439" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="14973" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="7981" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="7955" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="7956" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="7957" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="7984" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="7985" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="7986" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="7988" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="7987" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="7989" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="7958" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="7959" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="7960" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="7961" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="7962" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="7963" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="7964" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="7965" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="7966" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="7967" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="7968" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="7969" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="7970" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="7971" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="7972" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="7973" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="7974" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="7975" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="7976" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="7978" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="7979" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="14974" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18440" agemax="-1" agemin="17" name="Classe S16-Senior" handicap="16" />
                <AGEGROUP agegroupid="18441" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="8925" agemax="-1" agemin="17" name="Classe S17-Senior" handicap="17" />
                <AGEGROUP agegroupid="7982" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="7983" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="11114" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="8926" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="14975" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2448" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="650" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15310" agemax="-1" agemin="-1" name="Classe S14-Absolutos" />
                <AGEGROUP agegroupid="15314" agemax="-1" agemin="-1" name="Classe S21 (SDown)-Absolutos" />
                <AGEGROUP agegroupid="15320" agemax="-1" agemin="-1" name="34 Pontos-Abs" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2023-12-02" daytime="15:30" endtime="18:07" name="1ª Jornada - 2ª Sessão" number="2" warmupfrom="14:00" warmupuntil="15:15" maxentriesathlete="2">
          <EVENTS>
            <EVENT eventid="1143" daytime="15:30" gender="F" number="16" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="7888" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="7901" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="14976" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18152" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="7905" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="7889" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="7890" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="7891" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="7892" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="20872" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="20873" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="7908" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="7909" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="7923" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="7922" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="7910" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="7911" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="7921" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="7912" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="7920" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="7913" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="7919" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="7914" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="7918" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="7915" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="7917" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="7916" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="7899" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="7900" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="7902" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="7903" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="9886" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="14977" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18153" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18154" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="7906" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="7907" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="11115" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="7904" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="14978" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1151" gender="M" number="17" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="20874" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="20875" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="20876" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="20877" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="20878" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="20879" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="20880" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="20881" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="20882" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="20883" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="20884" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="20885" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="20886" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="20887" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="20888" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="20889" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="20890" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="20891" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="20892" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="20893" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="20894" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="20895" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="20896" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="20897" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="20898" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="20899" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="20900" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="20901" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="20902" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="20903" agemax="16" agemin="8" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="20904" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="20905" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="20906" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="20907" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="20908" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="20909" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="20910" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="20911" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="20912" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="20913" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5886" gender="F" number="18" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18524" agemax="-1" agemin="10" name="Classe S14-Absoluto" handicap="14" />
                <AGEGROUP agegroupid="7692" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absoluto" handicap="15" />
                <AGEGROUP agegroupid="7689" agemax="-1" agemin="10" name="Classe S17-Absoluto" handicap="17" />
                <AGEGROUP agegroupid="7695" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absoluto" handicap="21" />
                <AGEGROUP agegroupid="7690" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18526" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18525" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="7691" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="7693" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="7694" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="7696" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="7697" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="5901" gender="M" number="19" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18527" agemax="-1" agemin="10" name="Classe S14-Absoluto" handicap="14" />
                <AGEGROUP agegroupid="18528" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absoluto" handicap="15" />
                <AGEGROUP agegroupid="18529" agemax="-1" agemin="10" name="Classe S17-Absoluto" handicap="17" />
                <AGEGROUP agegroupid="18530" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absoluto" handicap="21" />
                <AGEGROUP agegroupid="18531" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18532" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18533" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18534" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18535" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18536" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18537" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18538" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1070" gender="F" number="20" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18380" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,14" />
                <AGEGROUP agegroupid="18381" agemax="-1" agemin="8" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18382" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18383" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="18384" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="18385" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="18386" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="18387" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="18388" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="18389" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="18390" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="18391" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="18392" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="18393" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="18394" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="18395" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18396" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18397" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18398" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18399" agemax="-1" agemin="-1" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18400" agemax="-1" agemin="-1" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18401" agemax="-1" agemin="-1" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18402" agemax="-1" agemin="-1" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18403" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18404" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18405" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1058" gender="M" number="21" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="24576" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="24577" agemax="-1" agemin="8" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="24578" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="24579" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="24580" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="24581" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="24582" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="24583" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="24584" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="24585" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="24586" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="24587" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="24588" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="24589" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="24590" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="24591" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="24592" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="24593" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="24594" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="24595" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="24596" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="24597" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="24598" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="24599" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="24600" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="24601" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="24602" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="24603" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="24604" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="24605" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="24606" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="24607" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="24608" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="24609" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="24610" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="24611" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="24612" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="24613" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="24614" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="24615" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="24616" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="24617" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="24618" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="24619" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1168" gender="F" number="22" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="150" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12264" agemax="-1" agemin="10" name="Classe SM1-SM4-Absolutos" handicap="1,2,3,4" />
                <AGEGROUP agegroupid="12265" agemax="16" agemin="10" name="Classe SM1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="12266" agemax="-1" agemin="17" name="Classe SM1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="12267" agemax="16" agemin="10" name="Classe SM2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="12268" agemax="-1" agemin="17" name="Classe SM2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="12269" agemax="16" agemin="10" name="Classe SM3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="12270" agemax="-1" agemin="17" name="Classe SM3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="12271" agemax="16" agemin="10" name="Classe SM4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="12272" agemax="-1" agemin="17" name="Classe SM4-Seniores" handicap="4" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1159" gender="M" number="23" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="150" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2703" agemax="-1" agemin="10" name="Classe SM1-SM4-Absolutos" handicap="1,2,3,4" />
                <AGEGROUP agegroupid="8098" agemax="16" agemin="10" name="Classe SM1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="2699" agemax="-1" agemin="17" name="Classe SM1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="8100" agemax="16" agemin="10" name="Classe SM2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="2700" agemax="-1" agemin="17" name="Classe SM2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="2701" agemax="16" agemin="10" name="Classe SM3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="8101" agemax="-1" agemin="17" name="Classe SM3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="8102" agemax="16" agemin="10" name="Classe SM4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="2702" agemax="-1" agemin="17" name="Classe SM4-Seniores" handicap="4" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1191" gender="F" number="24" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18341" agemax="-1" agemin="10" name="Classe SM5-SM14-Absolutos" handicap="5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="18342" agemax="-1" agemin="10" name="Classe SM15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18343" agemax="-1" agemin="-1" name="Classe SM16-Absolutos" />
                <AGEGROUP agegroupid="18344" agemax="-1" agemin="-1" name="Classe SM17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="18345" agemax="-1" agemin="10" name="Classe SM21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="18346" agemax="16" agemin="10" name="Classe SM5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="18347" agemax="-1" agemin="17" name="Classe SM5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="18348" agemax="16" agemin="10" name="Classe SM6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="18349" agemax="-1" agemin="17" name="Classe SM6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="18350" agemax="16" agemin="10" name="Classe SM7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="18351" agemax="-1" agemin="17" name="Classe SM7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="18352" agemax="16" agemin="10" name="Classe SM8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="18353" agemax="-1" agemin="17" name="Classe SM8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="18354" agemax="17" agemin="10" name="Classe SM9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="18355" agemax="-1" agemin="17" name="Classe SM9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="18356" agemax="16" agemin="10" name="Classe SM10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="18357" agemax="-1" agemin="17" name="Classe SM10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="18358" agemax="16" agemin="10" name="Classe SM11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="18359" agemax="-1" agemin="17" name="Classe SM11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="18360" agemax="16" agemin="10" name="Classe SM12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="18361" agemax="-1" agemin="17" name="Classe SM12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="18362" agemax="16" agemin="10" name="Classe SM13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="18363" agemax="-1" agemin="17" name="Classe SM13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="18364" agemax="16" agemin="10" name="Classe SM14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18365" agemax="-1" agemin="17" name="Classe SM14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18366" agemax="16" agemin="10" name="Classe SM15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18367" agemax="-1" agemin="17" name="Classe SM15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18368" agemax="-1" agemin="-1" name="Classe SM16-Esperanças" />
                <AGEGROUP agegroupid="18369" agemax="-1" agemin="-1" name="Classe SM16-Seniores" />
                <AGEGROUP agegroupid="18370" agemax="-1" agemin="-1" name="Classe SM17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18371" agemax="-1" agemin="-1" name="Classe SM17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18372" agemax="16" agemin="10" name="Classe SM21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18373" agemax="-1" agemin="17" name="Classe SM21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18374" agemax="-1" agemin="-1" name="Classe SM110" handicap="110" />
                <AGEGROUP agegroupid="18375" agemax="-1" agemin="-1" name="Classe SM113" handicap="113" />
                <AGEGROUP agegroupid="18376" agemax="-1" agemin="-1" name="Classe SM114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1173" gender="M" number="25" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8126" agemax="-1" agemin="10" name="Classe SM5-SM14-Absolutos" handicap="5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="8122" agemax="-1" agemin="10" name="Classe SM15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18338" agemax="-1" agemin="-1" name="Classe SM16-Absolutos" />
                <AGEGROUP agegroupid="14991" agemax="-1" agemin="-1" name="Classe SM17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="8123" agemax="-1" agemin="10" name="Classe SM21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="8112" agemax="16" agemin="10" name="Classe SM5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="1189" agemax="-1" agemin="17" name="Classe SM5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="8113" agemax="16" agemin="10" name="Classe SM6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="1174" agemax="-1" agemin="17" name="Classe SM6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="8114" agemax="16" agemin="10" name="Classe SM7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="1175" agemax="-1" agemin="17" name="Classe SM7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="8115" agemax="16" agemin="10" name="Classe SM8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="1176" agemax="-1" agemin="17" name="Classe SM8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="8116" agemax="17" agemin="10" name="Classe SM9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="1177" agemax="-1" agemin="17" name="Classe SM9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="8117" agemax="16" agemin="10" name="Classe SM10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="1931" agemax="-1" agemin="17" name="Classe SM10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="8118" agemax="16" agemin="10" name="Classe SM11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="1932" agemax="-1" agemin="17" name="Classe SM11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="8119" agemax="16" agemin="10" name="Classe SM12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="4024" agemax="-1" agemin="17" name="Classe SM12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="8120" agemax="16" agemin="10" name="Classe SM13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="1178" agemax="-1" agemin="17" name="Classe SM13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="8121" agemax="16" agemin="10" name="Classe SM14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="1179" agemax="-1" agemin="17" name="Classe SM14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="8125" agemax="16" agemin="10" name="Classe SM15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="6084" agemax="-1" agemin="17" name="Classe SM15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="14990" agemax="-1" agemin="-1" name="Classe SM16-Esperanças" />
                <AGEGROUP agegroupid="6345" agemax="-1" agemin="-1" name="Classe SM16-Seniores" />
                <AGEGROUP agegroupid="18339" agemax="-1" agemin="-1" name="Classe SM17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18340" agemax="-1" agemin="-1" name="Classe SM17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="1953" agemax="16" agemin="10" name="Classe SM21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="8124" agemax="-1" agemin="17" name="Classe SM21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="3267" agemax="-1" agemin="-1" name="Classe SM110" handicap="110" />
                <AGEGROUP agegroupid="6346" agemax="-1" agemin="-1" name="Classe SM113" handicap="113" />
                <AGEGROUP agegroupid="14992" agemax="-1" agemin="-1" name="Classe SM114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1215" gender="F" number="26" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8209" agemax="-1" agemin="10" name="Classe SB1-SB14-Absolutos" handicap="1,2,3,4,5,6,7,14" />
                <AGEGROUP agegroupid="8238" agemax="-1" agemin="10" name="Classe SB15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="15000" agemax="-1" agemin="-1" name="Classe SB16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="19518" agemax="-1" agemin="-1" name="Classe SB17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="8242" agemax="-1" agemin="10" name="Classe SB21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="8210" agemax="-1" agemin="17" name="Classe SB1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="8211" agemax="16" agemin="10" name="Classe SB1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="8212" agemax="16" agemin="10" name="Classe SB2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="8213" agemax="-1" agemin="17" name="Classe SB2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="8214" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="8215" agemax="-1" agemin="17" name="Classe SB3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="8216" agemax="16" agemin="10" name="Classe SB4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="8217" agemax="-1" agemin="17" name="Classe SB14-Seniores" handicap="4" />
                <AGEGROUP agegroupid="8218" agemax="16" agemin="10" name="Classe SB15-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="8219" agemax="-1" agemin="17" name="Classe SB15-Seniores" handicap="5" />
                <AGEGROUP agegroupid="8220" agemax="16" agemin="10" name="Classe SB16-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="8221" agemax="-1" agemin="17" name="Classe SB16-Seniores" handicap="6" />
                <AGEGROUP agegroupid="8222" agemax="16" agemin="10" name="Classe SB17-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="8223" agemax="-1" agemin="17" name="Classe SB17-Seniores" handicap="7" />
                <AGEGROUP agegroupid="8243" agemax="16" agemin="10" name="Classe SB21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="8244" agemax="-1" agemin="17" name="Classe SB21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="8241" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23338" gender="M" number="27" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23339" agemax="-1" agemin="10" name="Classe SB1-SB14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="23340" agemax="-1" agemin="10" name="Classe SB15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="23341" agemax="-1" agemin="-1" name="Classe SB16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="23342" agemax="-1" agemin="-1" name="Classe SB17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="23343" agemax="-1" agemin="10" name="Classe SB21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="23344" agemax="-1" agemin="17" name="Classe SB1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="23345" agemax="16" agemin="10" name="Classe SB1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="23346" agemax="16" agemin="10" name="Classe SB2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="23347" agemax="-1" agemin="17" name="Classe SB2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="23348" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="23349" agemax="-1" agemin="17" name="Classe SB3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="23350" agemax="16" agemin="10" name="Classe SB4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="23351" agemax="-1" agemin="17" name="Classe SB14-Seniores" handicap="4" />
                <AGEGROUP agegroupid="23352" agemax="16" agemin="10" name="Classe SB15-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="23353" agemax="-1" agemin="17" name="Classe SB15-Seniores" handicap="5" />
                <AGEGROUP agegroupid="23354" agemax="16" agemin="10" name="Classe SB16-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="23355" agemax="-1" agemin="17" name="Classe SB16-Seniores" handicap="6" />
                <AGEGROUP agegroupid="23356" agemax="16" agemin="10" name="Classe SB17-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="23357" agemax="-1" agemin="17" name="Classe SB17-Seniores" handicap="7" />
                <AGEGROUP agegroupid="23358" agemax="16" agemin="10" name="Classe SB21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="23359" agemax="-1" agemin="17" name="Classe SB21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="23360" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="24620" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1225" gender="F" number="28" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12321" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,14" />
                <AGEGROUP agegroupid="12338" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="19521" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="15002" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="12342" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="12322" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="12323" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="12324" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="12325" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="12326" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="12327" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="12328" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="12329" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="12331" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="12330" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="12332" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="12333" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="12334" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="12335" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="12336" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="12337" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="12339" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="12340" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="15003" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="19522" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="19523" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="12341" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="12343" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="12344" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="12345" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="12346" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="23378" gender="M" number="29" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="23379" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,14" />
                <AGEGROUP agegroupid="23380" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="23381" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="23382" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="23383" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="23384" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="23385" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="23386" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="23387" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="23388" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="23389" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="23390" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="23391" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="23392" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="23393" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="23394" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="23395" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="23396" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="23397" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="23398" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="23399" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="23400" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="23401" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="23402" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="23403" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="23404" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="23405" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="23406" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="23407" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="23408" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="23409" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1134" gender="F" number="30" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="12347" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="12376" agemax="-1" agemin="10" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18276" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="15004" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="12380" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="12348" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="12349" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="12350" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="12351" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="12352" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="12353" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="12354" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="12355" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="12356" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="12357" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="12358" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="12359" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="12360" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="12361" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="12362" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="12363" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="12364" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="12365" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="12366" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="12367" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="12368" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="12369" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="12370" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="12371" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="12372" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="12373" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="12374" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="12375" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="12377" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="12378" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18277" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18278" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="15005" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="12379" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="12381" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="12382" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="12383" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="12384" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="12385" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1138" gender="M" number="31" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="18279" agemax="-1" agemin="10" name="Classe S1-S14-Absolutos" handicap="1,2,3,4,5,6,7,8,9,10,11,12,13,14" />
                <AGEGROUP agegroupid="18280" agemax="-1" agemin="8" name="Classe S15 (Auditiva)-Absolutos" handicap="15" />
                <AGEGROUP agegroupid="18281" agemax="-1" agemin="-1" name="Classe S16-Absolutos" handicap="16" />
                <AGEGROUP agegroupid="18282" agemax="-1" agemin="-1" name="Classe S17-Absolutos" handicap="17" />
                <AGEGROUP agegroupid="18283" agemax="-1" agemin="10" name="Classe S21 (SDown)-Absolutos" handicap="21" />
                <AGEGROUP agegroupid="18284" agemax="16" agemin="10" name="Classe S1-Esperanças" handicap="1" />
                <AGEGROUP agegroupid="18285" agemax="-1" agemin="17" name="Classe S1-Seniores" handicap="1" />
                <AGEGROUP agegroupid="18286" agemax="16" agemin="10" name="Classe S2-Esperanças" handicap="2" />
                <AGEGROUP agegroupid="18287" agemax="-1" agemin="17" name="Classe S2-Seniores" handicap="2" />
                <AGEGROUP agegroupid="18288" agemax="16" agemin="10" name="Classe S3-Esperanças" handicap="3" />
                <AGEGROUP agegroupid="18289" agemax="-1" agemin="17" name="Classe S3-Seniores" handicap="3" />
                <AGEGROUP agegroupid="18290" agemax="16" agemin="10" name="Classe S4-Esperanças" handicap="4" />
                <AGEGROUP agegroupid="18291" agemax="-1" agemin="17" name="Classe S4-Seniores" handicap="4" />
                <AGEGROUP agegroupid="18292" agemax="16" agemin="10" name="Classe S5-Esperanças" handicap="5" />
                <AGEGROUP agegroupid="18293" agemax="-1" agemin="17" name="Classe S5-Seniores" handicap="5" />
                <AGEGROUP agegroupid="18294" agemax="16" agemin="10" name="Classe S6-Esperanças" handicap="6" />
                <AGEGROUP agegroupid="18295" agemax="-1" agemin="17" name="Classe S6-Seniores" handicap="6" />
                <AGEGROUP agegroupid="18296" agemax="16" agemin="10" name="Classe S7-Esperanças" handicap="7" />
                <AGEGROUP agegroupid="18297" agemax="-1" agemin="17" name="Classe S7-Seniores" handicap="7" />
                <AGEGROUP agegroupid="18298" agemax="16" agemin="10" name="Classe S8-Esperanças" handicap="8" />
                <AGEGROUP agegroupid="18299" agemax="-1" agemin="17" name="Classe S8-Seniores" handicap="8" />
                <AGEGROUP agegroupid="18300" agemax="16" agemin="10" name="Classe S9-Esperanças" handicap="9" />
                <AGEGROUP agegroupid="18301" agemax="-1" agemin="17" name="Classe S9-Seniores" handicap="9" />
                <AGEGROUP agegroupid="18302" agemax="16" agemin="10" name="Classe S10-Esperanças" handicap="10" />
                <AGEGROUP agegroupid="18303" agemax="-1" agemin="17" name="Classe S10-Seniores" handicap="10" />
                <AGEGROUP agegroupid="18304" agemax="16" agemin="10" name="Classe S11-Esperanças" handicap="11" />
                <AGEGROUP agegroupid="18305" agemax="-1" agemin="17" name="Classe S11-Seniores" handicap="11" />
                <AGEGROUP agegroupid="18306" agemax="16" agemin="10" name="Classe S12-Esperanças" handicap="12" />
                <AGEGROUP agegroupid="18307" agemax="-1" agemin="17" name="Classe S12-Seniores" handicap="12" />
                <AGEGROUP agegroupid="18308" agemax="16" agemin="10" name="Classe S13-Esperanças" handicap="13" />
                <AGEGROUP agegroupid="18309" agemax="-1" agemin="17" name="Classe S13-Seniores" handicap="13" />
                <AGEGROUP agegroupid="18310" agemax="16" agemin="10" name="Classe S14-Esperanças" handicap="14" />
                <AGEGROUP agegroupid="18311" agemax="-1" agemin="17" name="Classe S14-Seniores" handicap="14" />
                <AGEGROUP agegroupid="18312" agemax="16" agemin="10" name="Classe S15 (Auditiva)-Esperanças" handicap="15" />
                <AGEGROUP agegroupid="18313" agemax="-1" agemin="17" name="Classe S15 (Auditiva)-Seniores" handicap="15" />
                <AGEGROUP agegroupid="18314" agemax="16" agemin="10" name="Classe S16-Esperanças" handicap="16" />
                <AGEGROUP agegroupid="18315" agemax="-1" agemin="17" name="Classe S16-Seniores" handicap="16" />
                <AGEGROUP agegroupid="18316" agemax="16" agemin="10" name="Classe S17-Esperanças" handicap="17" />
                <AGEGROUP agegroupid="18317" agemax="-1" agemin="17" name="Classe S17-Seniores" handicap="17" />
                <AGEGROUP agegroupid="18318" agemax="16" agemin="10" name="Classe S21 (SDown)-Esperanças" handicap="21" />
                <AGEGROUP agegroupid="18319" agemax="-1" agemin="17" name="Classe S21 (SDown)-Seniores" handicap="21" />
                <AGEGROUP agegroupid="18320" agemax="-1" agemin="-1" name="Classe S110" handicap="110" />
                <AGEGROUP agegroupid="18321" agemax="-1" agemin="-1" name="Classe S113" handicap="113" />
                <AGEGROUP agegroupid="18322" agemax="-1" agemin="-1" name="Classe S114" handicap="114" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="2496" number="32" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="650" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="15338" agemax="-1" agemin="-1" name="Classe S14-Absolutos" />
                <AGEGROUP agegroupid="15339" agemax="-1" agemin="-1" name="Classe S21 (SDown)-Absolutos" />
                <AGEGROUP agegroupid="15340" agemax="-1" agemin="-1" name="34 Pontos-Abs" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
    </MEET>
  </MEETS>
</LENEX>
