<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Team Manager 10" registration="Clube Nautico Academico" version="10.75980">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET name="Campeonato Interdistrital de Juvenis, Juniores e Seniores PL" number="20" city="Coimbra" nation="POR" deadline="2023-07-05" course="LCM">
      <POOL name="Centro Olimpico de Piscinas" />
      <AGEDATE value="2023-07-14" type="POR" />
      <QUALIFY from="2022-07-11" until="2023-07-03" />
      <SESSIONS>
        <SESSION number="1" date="2023-07-14" daytime="16:30">
          <EVENTS>
            <EVENT number="1" gender="M" eventid="10" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="2" gender="F" eventid="20" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="3" gender="M" eventid="30" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="4" gender="F" eventid="40" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2023-07-15" daytime="09:00">
          <EVENTS>
            <EVENT number="5" gender="M" eventid="50" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="6" gender="F" eventid="60" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="7" gender="M" eventid="70" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="8" gender="F" eventid="80" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="9" gender="M" eventid="90" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="10" gender="F" eventid="100" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="11" gender="M" eventid="110" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="12" gender="F" eventid="120" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="13" gender="M" eventid="130" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="14" gender="F" eventid="140" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="3" date="2023-07-15" daytime="16:00">
          <EVENTS>
            <EVENT number="15" eventid="150" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemin="14" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="16" gender="F" eventid="160" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="17" gender="M" eventid="170" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="18" gender="F" eventid="180" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="19" gender="M" eventid="190" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="20" gender="F" eventid="200" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="21" gender="M" eventid="210" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="22" gender="F" eventid="220" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="23" gender="M" eventid="230" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="24" gender="M" eventid="240" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="25" gender="F" eventid="250" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="4" date="2023-07-16" daytime="09:00">
          <EVENTS>
            <EVENT number="26" gender="F" eventid="260" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="27" gender="M" eventid="270" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="28" gender="F" eventid="280" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="29" gender="M" eventid="290" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="-1" />
                <AGEGROUP agegroupid="2" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="30" gender="F" eventid="300" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="31" gender="M" eventid="310" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="32" gender="F" eventid="320" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="33" gender="M" eventid="330" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="34" gender="F" eventid="340" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="35" gender="M" eventid="350" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="36" eventid="360" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" agemin="14" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="5" date="2023-07-16" daytime="16:00">
          <EVENTS>
            <EVENT number="37" gender="M" eventid="370" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="38" gender="F" eventid="380" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="39" gender="M" eventid="390" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="40" gender="F" eventid="400" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="41" gender="M" eventid="410" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="42" gender="F" eventid="420" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="43" gender="M" eventid="430" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="2" gender="M" agemin="16" agemax="16" />
                <AGEGROUP agegroupid="3" gender="M" agemin="17" agemax="18" />
                <AGEGROUP agegroupid="4" gender="M" agemin="19" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="44" gender="F" eventid="440" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE value="260" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="14" />
                <AGEGROUP agegroupid="2" gender="F" agemin="15" agemax="15" />
                <AGEGROUP agegroupid="3" gender="F" agemin="16" agemax="17" />
                <AGEGROUP agegroupid="4" gender="F" agemin="18" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="45" gender="M" eventid="450" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="M" agemin="15" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
            <EVENT number="46" gender="F" eventid="460" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE value="750" currency="EUR" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1" gender="F" agemin="14" agemax="-1" />
              </AGEGROUPS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB clubid="6" name="Clube Náutico Académico de Coimbra" shortname="CNAC" code="CNAC" nation="POR" region="ANC">
          <ATHLETES>
            <ATHLETE athleteid="3933" lastname="Aguilar" firstname="Marta Andre" gender="F" license="132766" birthdate="2007-03-14">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:18:27.74">
                  <MEETINFO course="LCM" date="2023-02-12" city="Lisboa" nation="POR" name="ARENA LISBON INTERNATIONAL MEETING 2023" />
                </ENTRY>
                <ENTRY eventid="100" entrytime="00:01:03.97">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="220" entrytime="00:02:16.78">
                  <MEETINFO course="LCM" date="2023-02-11" city="Lisboa" nation="POR" name="ARENA LISBON INTERNATIONAL MEETING 2023" />
                </ENTRY>
                <ENTRY eventid="280" entrytime="00:09:39.35">
                  <MEETINFO course="LCM" date="2023-05-27" city="Coimbra" nation="POR" name="XV Meeting Cidade de Coimbra / XXXIV TQueima das Fitas" />
                </ENTRY>
                <ENTRY eventid="420" entrytime="00:04:42.21">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="300" entrytime="00:00:30.04">
                  <MEETINFO course="LCM" date="2023-04-29" city="Coimbra" nation="POR" name="XXXVII Torneio de Natação do CNAC- Shigeo Tsukagoshi" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4373" lastname="Almeida" firstname="Joao Neves" gender="M" license="129566" birthdate="2005-01-20">
              <ENTRIES>
                <ENTRY eventid="70" entrytime="00:09:17.38">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="170" entrytime="00:01:03.75">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="330" entrytime="00:02:16.27">
                  <MEETINFO course="LCM" date="2023-05-28" city="Coimbra" nation="POR" name="XV Meeting Cidade de Coimbra / XXXIV TQueima das Fitas" />
                </ENTRY>
                <ENTRY eventid="410" entrytime="00:04:29.26">
                  <MEETINFO course="LCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="264" lastname="Bastos" firstname="Lucas Pereira" gender="M" license="117492" birthdate="2000-08-03">
              <ENTRIES>
                <ENTRY eventid="110" entrytime="00:02:17.20">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="230" entrytime="00:01:55.24">
                  <MEETINFO course="LCM" date="2023-04-02" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="290" entrytime="00:04:32.11">
                  <MEETINFO course="LCM" date="2022-07-28" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="410" entrytime="00:04:04.81">
                  <MEETINFO course="LCM" date="2023-04-01" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="430" entrytime="00:02:11.26">
                  <MEETINFO course="LCM" date="2023-04-01" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="350" entrytime="00:01:07.38">
                  <MEETINFO course="LCM" date="2023-04-06" city="Oeiras" nation="POR" name="Campeonato Nacional Clubes 1 Divisão" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="812" lastname="Bastos" firstname="Vasco Pereira" gender="M" license="119766" birthdate="2002-09-11">
              <ENTRIES>
                <ENTRY eventid="90" entrytime="00:00:54.05">
                  <MEETINFO course="LCM" date="2023-03-31" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="130" entrytime="00:00:31.45">
                  <MEETINFO course="LCM" date="2023-04-07" city="Oeiras" nation="POR" name="Campeonato Nacional Clubes 1 Divisão" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4731" lastname="Cortesao" firstname="Maria Manuel" gender="F" license="203972" birthdate="2008-10-17">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:19:22.04">
                  <MEETINFO course="LCM" date="2023-03-30" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="100" entrytime="00:01:05.38">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="220" entrytime="00:02:22.67">
                  <MEETINFO course="LCM" date="2023-02-11" city="Lisboa" nation="POR" name="ARENA LISBON INTERNATIONAL MEETING 2023" />
                </ENTRY>
                <ENTRY eventid="280" entrytime="00:10:12.21">
                  <MEETINFO course="LCM" date="2023-03-31" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="420" entrytime="00:05:00.81">
                  <MEETINFO course="LCM" date="2023-04-01" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4984" lastname="Cruz" firstname="Ana Margarida" gender="F" license="208419" sdmsid="0" birthdate="2009-11-10">
              <ENTRIES>
                <ENTRY eventid="140" entrytime="00:00:39.59">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="220" entrytime="00:02:26.78">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="300" entrytime="00:00:31.35">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="340" entrytime="00:01:33.31">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="420" entrytime="00:05:14.87">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4950" lastname="Cunha" firstname="Joaquim Antonio" gender="M" license="205507" birthdate="2008-07-25">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:18:25.84">
                  <MEETINFO course="LCM" date="2023-03-17" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="70" entrytime="00:09:55.81">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="230" entrytime="00:02:19.25">
                  <MEETINFO course="LCM" date="2023-04-29" city="Coimbra" nation="POR" name="XXXVII Torneio de Natação do CNAC- Shigeo Tsukagoshi" />
                </ENTRY>
                <ENTRY eventid="290" entrytime="00:05:31.47">
                  <MEETINFO course="SCM" date="2023-05-21" city="Cantanhede" nation="POR" name="Torneio Regional de Fundo Infantis e Juvenis" />
                </ENTRY>
                <ENTRY eventid="410" entrytime="00:04:54.10">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="2621" lastname="Diogo" firstname="Dinis Miranda" gender="M" license="129397" birthdate="2004-09-22">
              <ENTRIES>
                <ENTRY eventid="110" entrytime="00:02:24.18">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="190" entrytime="00:00:29.59">
                  <MEETINFO course="LCM" date="2023-01-22" city="Coimbra" nation="POR" name="Taça Velocidade" />
                </ENTRY>
                <ENTRY eventid="350" entrytime="00:01:16.27">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="370" entrytime="00:01:02.41">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="430" entrytime="00:02:15.23">
                  <MEETINFO course="LCM" date="2022-07-30" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4653" lastname="Diogo" firstname="Ines Miranda" gender="F" license="200416" birthdate="2007-10-16">
              <ENTRIES>
                <ENTRY eventid="120" entrytime="00:02:34.40">
                  <MEETINFO course="LCM" date="2022-12-17" city="Coimbra" nation="POR" name="2022 Coimbra Swimming OPEN" />
                </ENTRY>
                <ENTRY eventid="180" entrytime="00:00:34.37">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="220" entrytime="00:02:15.22">
                  <MEETINFO course="LCM" date="2023-02-11" city="Lisboa" nation="POR" name="ARENA LISBON INTERNATIONAL MEETING 2023" />
                </ENTRY>
                <ENTRY eventid="280" entrytime="00:09:49.97">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="380" entrytime="00:01:12.30">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="420" entrytime="00:04:44.46">
                  <MEETINFO course="LCM" date="2023-02-12" city="Lisboa" nation="POR" name="ARENA LISBON INTERNATIONAL MEETING 2023" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="5140" lastname="Domingues" firstname="Ana Beatriz" gender="F" license="216734" birthdate="2008-02-05">
              <ENTRIES>
                <ENTRY eventid="100" entrytime="00:01:09.27">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="180" entrytime="00:00:34.77">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="300" entrytime="00:00:31.23">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="400" entrytime="00:00:32.91">
                  <MEETINFO course="LCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4962" lastname="Fernandes" firstname="Laura Carvalho" gender="F" license="208551" birthdate="2008-12-15">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:20:15.55">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="80" entrytime="00:05:49.20">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="160" entrytime="00:01:14.72">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="320" entrytime="00:02:48.23">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="420" entrytime="00:05:03.92">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4377" lastname="Ferreira" firstname="Joao Rafael" gender="M" license="148624" birthdate="2006-07-18">
              <ENTRIES>
                <ENTRY eventid="90" entrytime="00:00:57.90">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="230" entrytime="00:02:07.63">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="310" entrytime="00:00:26.17">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="3938" lastname="Ferreira" firstname="Maria Neto" gender="F" license="131467" birthdate="2006-08-24">
              <ENTRIES>
                <ENTRY eventid="40" entrytime="00:19:12.38">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="160" entrytime="00:01:07.92">
                  <MEETINFO course="LCM" date="2022-12-17" city="Coimbra" nation="POR" name="2022 Coimbra Swimming OPEN" />
                </ENTRY>
                <ENTRY eventid="220" entrytime="00:02:12.52">
                  <MEETINFO course="LCM" date="2022-07-28" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="320" entrytime="00:02:27.54">
                  <MEETINFO course="LCM" date="2023-03-30" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="420" entrytime="00:04:38.96">
                  <MEETINFO course="LCM" date="2023-04-01" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4619" lastname="Gaspar" firstname="Beatriz Andre" gender="F" license="132656" birthdate="2006-12-01">
              <ENTRIES>
                <ENTRY eventid="140" entrytime="00:00:37.99">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="200" entrytime="00:02:44.78">
                  <MEETINFO course="LCM" date="2022-07-29" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="340" entrytime="00:01:17.72">
                  <MEETINFO course="LCM" date="2022-07-27" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="3942" lastname="Jesus" firstname="David Duarte" gender="M" license="131743" birthdate="2007-05-11">
              <ENTRIES>
                <ENTRY eventid="90" entrytime="00:00:59.47">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="230" entrytime="00:02:10.44">
                  <MEETINFO course="LCM" />
                </ENTRY>
                <ENTRY eventid="310" entrytime="00:00:26.89">
                  <MEETINFO course="LCM" date="2023-01-22" city="Coimbra" nation="POR" name="Taça Velocidade" />
                </ENTRY>
                <ENTRY eventid="410" entrytime="00:04:31.14">
                  <MEETINFO course="LCM" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4381" lastname="Mano" firstname="Leonor Mil" gender="F" license="202991" birthdate="2007-12-13">
              <ENTRIES>
                <ENTRY eventid="100" entrytime="00:00:59.71">
                  <MEETINFO course="LCM" date="2023-03-31" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="160" entrytime="00:01:09.01">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="220" entrytime="00:02:11.42">
                  <MEETINFO course="LCM" date="2023-05-27" city="Coimbra" nation="POR" name="XV Meeting Cidade de Coimbra / XXXIV TQueima das Fitas" />
                </ENTRY>
                <ENTRY eventid="300" entrytime="00:00:27.52">
                  <MEETINFO course="LCM" date="2023-03-30" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="400" entrytime="00:00:29.52">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4383" lastname="Oliveira" firstname="Carlos Miguel" gender="M" license="202983" birthdate="2006-01-09" />
            <ATHLETE athleteid="4961" lastname="Oliveira" firstname="Marco Dimitar" gender="M" license="209588" birthdate="2007-02-01">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:17:30.52">
                  <MEETINFO course="LCM" date="2023-03-17" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="70" entrytime="00:09:12.29">
                  <MEETINFO course="LCM" date="2023-03-31" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="230" entrytime="00:02:09.72">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="410" entrytime="00:04:34.04">
                  <MEETINFO course="LCM" date="2023-04-01" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4387" lastname="Pereira" firstname="Tomas Veiga" gender="M" license="137055" birthdate="2006-07-06">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:17:33.66">
                  <MEETINFO course="LCM" date="2022-07-27" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="70" entrytime="00:09:13.35">
                  <MEETINFO course="LCM" date="2022-07-30" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="170" entrytime="00:01:04.54">
                  <MEETINFO course="LCM" date="2023-04-29" city="Coimbra" nation="POR" name="XXXVII Torneio de Natação do CNAC- Shigeo Tsukagoshi" />
                </ENTRY>
                <ENTRY eventid="330" entrytime="00:02:20.97">
                  <MEETINFO course="LCM" date="2023-04-06" city="Oeiras" nation="POR" name="Campeonato Nacional Clubes 1 Divisão" />
                </ENTRY>
                <ENTRY eventid="410" entrytime="00:04:27.00">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="3721" lastname="Reis" firstname="Rodrigo Miguel" gender="M" license="129842" birthdate="2004-05-28">
              <ENTRIES>
                <ENTRY eventid="90" entrytime="00:00:53.32">
                  <MEETINFO course="LCM" date="2023-03-31" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="170" entrytime="00:00:57.95">
                  <MEETINFO course="LCM" date="2022-07-29" city="Oeiras" nation="POR" name="Campeonatos Nacionais Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="310" entrytime="00:00:24.32">
                  <MEETINFO course="LCM" date="2023-03-30" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="390" entrytime="00:00:25.98">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="5143" lastname="Silveira" firstname="Gabriela Luca" gender="F" license="219176" birthdate="2009-03-25" />
            <ATHLETE athleteid="4391" lastname="Sousa" firstname="Guilherme Simoes" gender="M" license="202988" birthdate="2008-11-26">
              <ENTRIES>
                <ENTRY eventid="30" entrytime="00:17:41.76">
                  <MEETINFO course="LCM" date="2023-03-30" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="70" entrytime="00:09:22.19">
                  <MEETINFO course="LCM" date="2023-03-31" city="Funchal" nation="POR" name="Campeonato Nacional Juvenis e Absolutos de Portugal OPEN" />
                </ENTRY>
                <ENTRY eventid="230" entrytime="00:02:10.93">
                  <MEETINFO course="LCM" date="2023-03-18" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
                <ENTRY eventid="350" entrytime="00:01:19.70">
                  <MEETINFO course="LCM" date="2023-06-24" city="Coimbra" nation="POR" name="Taça ANC" />
                </ENTRY>
                <ENTRY eventid="410" entrytime="00:04:33.90">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="1428" lastname="Travassos" firstname="Rodrigo Alexandre" gender="M" license="126187" birthdate="2002-08-06">
              <ENTRIES>
                <ENTRY eventid="90" entrytime="00:00:54.15">
                  <MEETINFO course="LCM" date="2023-04-07" city="Oeiras" nation="POR" name="Campeonato Nacional Clubes 1 Divisão" />
                </ENTRY>
                <ENTRY eventid="170" entrytime="00:00:59.86">
                  <MEETINFO course="LCM" date="2023-04-29" city="Coimbra" nation="POR" name="XXXVII Torneio de Natação do CNAC- Shigeo Tsukagoshi" />
                </ENTRY>
                <ENTRY eventid="310" entrytime="00:00:25.39">
                  <MEETINFO course="LCM" date="2023-04-29" city="Coimbra" nation="POR" name="XXXVII Torneio de Natação do CNAC- Shigeo Tsukagoshi" />
                </ENTRY>
                <ENTRY eventid="390" entrytime="00:00:27.17">
                  <MEETINFO course="LCM" date="2022-12-17" city="Coimbra" nation="POR" name="2022 Coimbra Swimming OPEN" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
            <ATHLETE athleteid="4618" lastname="Varela" firstname="Joana Filipa" gender="F" license="133977" birthdate="2006-10-07">
              <ENTRIES>
                <ENTRY eventid="180" entrytime="00:00:36.09">
                  <MEETINFO course="LCM" date="2022-12-17" city="Coimbra" nation="POR" name="2022 Coimbra Swimming OPEN" />
                </ENTRY>
                <ENTRY eventid="300" entrytime="00:00:31.27">
                  <MEETINFO course="LCM" date="2023-04-29" city="Coimbra" nation="POR" name="XXXVII Torneio de Natação do CNAC- Shigeo Tsukagoshi" />
                </ENTRY>
                <ENTRY eventid="400" entrytime="00:00:32.21">
                  <MEETINFO course="LCM" date="2023-03-19" city="Coimbra" nation="POR" name="Campeonato Interdistrital Juvenis, Juniores e Absolutos PL" />
                </ENTRY>
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY relayid="1" number="1" gender="M" agetotalmin="-1" agetotalmax="-1" agemin="17" agemax="18">
              <ENTRIES>
                <ENTRY eventid="270" entrytime="00:02:06.71">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4377">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4383">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4373">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4387">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="10" entrytime="00:08:40.53">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4373">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4387">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4377">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4383">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="50" entrytime="00:01:50.88">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4373">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4383">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4387">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4377">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="240" entrytime="00:03:56.27">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4373">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4387">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4383">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4377">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY relayid="2" number="1" gender="M" agetotalmin="-1" agetotalmax="-1" agemin="15" agemax="-1">
              <ENTRIES>
                <ENTRY eventid="450" entrytime="00:04:30.49">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4377">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4383">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4373">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4387">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY relayid="3" number="2" gender="M" agetotalmin="-1" agetotalmax="-1" agemin="19" agemax="-1">
              <ENTRIES>
                <ENTRY eventid="10" entrytime="00:07:59.63">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="264">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="1428">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="812">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3721">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="50" entrytime="00:01:45.25">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="264">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="812">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="1428">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3721">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="270" entrytime="00:01:56.01">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="2621">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="264">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="1428">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3721">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="450" entrytime="00:04:09.20">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="264">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="812">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="1428">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3721">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="240" entrytime="00:03:40.55">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="1428">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="264">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="2621">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3721">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY relayid="4" number="1" gender="F" agetotalmin="-1" agetotalmax="-1" agemin="16" agemax="17">
              <ENTRIES>
                <ENTRY eventid="20" entrytime="00:08:59.94">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4381">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="3933">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4653">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3938">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="60" entrytime="00:01:57.93">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4653">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4381">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="3933">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3938">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="250" entrytime="00:04:11.41">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4381">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="3933">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4653">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3938">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="260" entrytime="00:02:13.35">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4653">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4619">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4381">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3938">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="460" entrytime="00:04:41.65">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4653">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4619">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="3938">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4381">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY relayid="5" number="1" gender="X" agetotalmin="-1" agetotalmax="-1" agemin="14" agemax="15">
              <ENTRIES>
                <ENTRY eventid="150" entrytime="00:05:34.13">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4950">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4391">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4984">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="5143">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="360" entrytime="00:04:45.29">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4391">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4950">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4984">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="5143">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY relayid="6" number="2" gender="X" agetotalmin="-1" agetotalmax="-1" agemin="15" agemax="16">
              <ENTRIES>
                <ENTRY eventid="360" entrytime="00:04:20.69">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="3942">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4731">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4961">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4962">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="150" entrytime="00:04:58.33">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="3942">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4731">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4962">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4961">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
            <RELAY relayid="7" number="2" gender="X" agetotalmin="-1" agetotalmax="-1" agemin="16" agemax="18">
              <ENTRIES>
                <ENTRY eventid="360" entrytime="00:04:02.20">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4373">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4381">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="4377">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="3938">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
                <ENTRY eventid="150" entrytime="00:04:37.37">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="4373">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="2" athleteid="4383">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="3" athleteid="3938">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                    <RELAYPOSITION number="4" athleteid="4381">
                      <MEETINFO course="LCM" qualificationtime="NT" />
                    </RELAYPOSITION>
                  </RELAYPOSITIONS>
                </ENTRY>
              </ENTRIES>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
